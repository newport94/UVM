module counter (
                input wire [7:0] data_in,
                output reg [7:0] q,
                input wire clk,
                input wire inc, // counter increment
                input wire ld,  // bypass counter when high
                input wire rst);
`protected

    MTI!#j='O;.{l25c=Qm=;p?_|^73!O>$+!GRi]3!{N9?{'$~si[aa7e=<]sG}#To}QO[IszB~r1o
    7MZY_k2}5!F|!ax[B37zr[O,v{Iu&QCJT{B;[Ok_H<ITT!e2E<r5\u'O<]^AaML-5\-<(KnH~{}?
    _9=3*>$+vO,=r_+<>[P=QI]PjeeT2<}Wv3@{*bdp]vn3a]-
`endprotected
endmodule // counter
